// Copyright (C) 2019-2022 The SymbiFlow Authors
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC

module BANK();
	parameter FASM_EXTRA = "INTERNAL_VREF";
	parameter NUMBER = 0;
	parameter INTERNAL_VREF = 600;
endmodule
