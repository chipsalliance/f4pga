module GTPE2_CHANNEL (
    (* iopad_external_pin *)
    output GTPTXN,
    (* iopad_external_pin *)
    output GTPTXP,
    (* iopad_external_pin *)
    input GTPRXN,
    (* iopad_external_pin *)
    input GTPRXP
);

endmodule
