module \$_DFF_P_ (
    D,
    Q,
    C
);
  input D;
  input C;
  output Q;
  dff _TECHMAP_REPLACE_ (
      .Q  (Q),
      .D  (D),
      .CLK(C)
  );
endmodule

