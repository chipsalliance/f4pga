// Copyright 2020-2022 F4PGA Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// SPDX-License-Identifier: Apache-2.0

module top (
    input wire clk0,
    input wire clk1,
    (* clkbuf_inhibit *)
    input wire clk2,
    (* clkbuf_inhibit *)
    input wire clk3,

    input  wire [3:0] d,
    output reg  [3:0] q
);

  always @(posedge clk0) q[0] <= d[0];
  always @(posedge clk1) q[1] <= d[1];
  always @(posedge clk2) q[2] <= d[2];
  always @(posedge clk3) q[3] <= d[3];

endmodule
