module BANK();
	parameter FASM_EXTRA = "INTERNAL_VREF";
	parameter NUMBER = 0;
	parameter INTERNAL_VREF = 600;
endmodule
