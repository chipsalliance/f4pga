// Copyright (C) 2020-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier:ISC

module GTPE2_CHANNEL (
    (* iopad_external_pin *)
    output GTPTXN,
    (* iopad_external_pin *)
    output GTPTXP,
    (* iopad_external_pin *)
    input  GTPRXN,
    (* iopad_external_pin *)
    input  GTPRXP
);

endmodule
